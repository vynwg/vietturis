module c

#flag -luv

#include <uv.h>
