module c

#flag linux -L /usr/lib/
#flag linux -luv

#include <uv.h>
